// hps.v

// Generated using ACDS version 13.0sp1 232 at 2015.08.02.15:38:39

`timescale 1 ps / 1 ps
module hps (
		input  wire        clk_clk,                //            clk.clk
		input  wire        reset_reset_n,          //          reset.reset_n
		output wire [12:0] memory_mem_a,           //         memory.mem_a
		output wire [2:0]  memory_mem_ba,          //               .mem_ba
		output wire        memory_mem_ck,          //               .mem_ck
		output wire        memory_mem_ck_n,        //               .mem_ck_n
		output wire        memory_mem_cke,         //               .mem_cke
		output wire        memory_mem_cs_n,        //               .mem_cs_n
		output wire        memory_mem_ras_n,       //               .mem_ras_n
		output wire        memory_mem_cas_n,       //               .mem_cas_n
		output wire        memory_mem_we_n,        //               .mem_we_n
		output wire        memory_mem_reset_n,     //               .mem_reset_n
		inout  wire [7:0]  memory_mem_dq,          //               .mem_dq
		inout  wire        memory_mem_dqs,         //               .mem_dqs
		inout  wire        memory_mem_dqs_n,       //               .mem_dqs_n
		output wire        memory_mem_odt,         //               .mem_odt
		output wire        memory_mem_dm,          //               .mem_dm
		input  wire        memory_oct_rzqin,       //               .oct_rzqin
		output wire [11:0] h2f_axi_master_awid,    // h2f_axi_master.awid
		output wire [29:0] h2f_axi_master_awaddr,  //               .awaddr
		output wire [3:0]  h2f_axi_master_awlen,   //               .awlen
		output wire [2:0]  h2f_axi_master_awsize,  //               .awsize
		output wire [1:0]  h2f_axi_master_awburst, //               .awburst
		output wire [1:0]  h2f_axi_master_awlock,  //               .awlock
		output wire [3:0]  h2f_axi_master_awcache, //               .awcache
		output wire [2:0]  h2f_axi_master_awprot,  //               .awprot
		output wire        h2f_axi_master_awvalid, //               .awvalid
		input  wire        h2f_axi_master_awready, //               .awready
		output wire [11:0] h2f_axi_master_wid,     //               .wid
		output wire [63:0] h2f_axi_master_wdata,   //               .wdata
		output wire [7:0]  h2f_axi_master_wstrb,   //               .wstrb
		output wire        h2f_axi_master_wlast,   //               .wlast
		output wire        h2f_axi_master_wvalid,  //               .wvalid
		input  wire        h2f_axi_master_wready,  //               .wready
		input  wire [11:0] h2f_axi_master_bid,     //               .bid
		input  wire [1:0]  h2f_axi_master_bresp,   //               .bresp
		input  wire        h2f_axi_master_bvalid,  //               .bvalid
		output wire        h2f_axi_master_bready,  //               .bready
		output wire [11:0] h2f_axi_master_arid,    //               .arid
		output wire [29:0] h2f_axi_master_araddr,  //               .araddr
		output wire [3:0]  h2f_axi_master_arlen,   //               .arlen
		output wire [2:0]  h2f_axi_master_arsize,  //               .arsize
		output wire [1:0]  h2f_axi_master_arburst, //               .arburst
		output wire [1:0]  h2f_axi_master_arlock,  //               .arlock
		output wire [3:0]  h2f_axi_master_arcache, //               .arcache
		output wire [2:0]  h2f_axi_master_arprot,  //               .arprot
		output wire        h2f_axi_master_arvalid, //               .arvalid
		input  wire        h2f_axi_master_arready, //               .arready
		input  wire [11:0] h2f_axi_master_rid,     //               .rid
		input  wire [63:0] h2f_axi_master_rdata,   //               .rdata
		input  wire [1:0]  h2f_axi_master_rresp,   //               .rresp
		input  wire        h2f_axi_master_rlast,   //               .rlast
		input  wire        h2f_axi_master_rvalid,  //               .rvalid
		output wire        h2f_axi_master_rready   //               .rready
	);

	hps_hps_0 #(
		.F2S_Width (2),
		.S2F_Width (2)
	) hps_0 (
		.h2f_mpu_eventi     (),                       //    h2f_mpu_events.eventi
		.h2f_mpu_evento     (),                       //                  .evento
		.h2f_mpu_standbywfe (),                       //                  .standbywfe
		.h2f_mpu_standbywfi (),                       //                  .standbywfi
		.mem_a              (memory_mem_a),           //            memory.mem_a
		.mem_ba             (memory_mem_ba),          //                  .mem_ba
		.mem_ck             (memory_mem_ck),          //                  .mem_ck
		.mem_ck_n           (memory_mem_ck_n),        //                  .mem_ck_n
		.mem_cke            (memory_mem_cke),         //                  .mem_cke
		.mem_cs_n           (memory_mem_cs_n),        //                  .mem_cs_n
		.mem_ras_n          (memory_mem_ras_n),       //                  .mem_ras_n
		.mem_cas_n          (memory_mem_cas_n),       //                  .mem_cas_n
		.mem_we_n           (memory_mem_we_n),        //                  .mem_we_n
		.mem_reset_n        (memory_mem_reset_n),     //                  .mem_reset_n
		.mem_dq             (memory_mem_dq),          //                  .mem_dq
		.mem_dqs            (memory_mem_dqs),         //                  .mem_dqs
		.mem_dqs_n          (memory_mem_dqs_n),       //                  .mem_dqs_n
		.mem_odt            (memory_mem_odt),         //                  .mem_odt
		.mem_dm             (memory_mem_dm),          //                  .mem_dm
		.oct_rzqin          (memory_oct_rzqin),       //                  .oct_rzqin
		.h2f_rst_n          (),                       //         h2f_reset.reset_n
		.h2f_axi_clk        (clk_clk),                //     h2f_axi_clock.clk
		.h2f_AWID           (h2f_axi_master_awid),    //    h2f_axi_master.awid
		.h2f_AWADDR         (h2f_axi_master_awaddr),  //                  .awaddr
		.h2f_AWLEN          (h2f_axi_master_awlen),   //                  .awlen
		.h2f_AWSIZE         (h2f_axi_master_awsize),  //                  .awsize
		.h2f_AWBURST        (h2f_axi_master_awburst), //                  .awburst
		.h2f_AWLOCK         (h2f_axi_master_awlock),  //                  .awlock
		.h2f_AWCACHE        (h2f_axi_master_awcache), //                  .awcache
		.h2f_AWPROT         (h2f_axi_master_awprot),  //                  .awprot
		.h2f_AWVALID        (h2f_axi_master_awvalid), //                  .awvalid
		.h2f_AWREADY        (h2f_axi_master_awready), //                  .awready
		.h2f_WID            (h2f_axi_master_wid),     //                  .wid
		.h2f_WDATA          (h2f_axi_master_wdata),   //                  .wdata
		.h2f_WSTRB          (h2f_axi_master_wstrb),   //                  .wstrb
		.h2f_WLAST          (h2f_axi_master_wlast),   //                  .wlast
		.h2f_WVALID         (h2f_axi_master_wvalid),  //                  .wvalid
		.h2f_WREADY         (h2f_axi_master_wready),  //                  .wready
		.h2f_BID            (h2f_axi_master_bid),     //                  .bid
		.h2f_BRESP          (h2f_axi_master_bresp),   //                  .bresp
		.h2f_BVALID         (h2f_axi_master_bvalid),  //                  .bvalid
		.h2f_BREADY         (h2f_axi_master_bready),  //                  .bready
		.h2f_ARID           (h2f_axi_master_arid),    //                  .arid
		.h2f_ARADDR         (h2f_axi_master_araddr),  //                  .araddr
		.h2f_ARLEN          (h2f_axi_master_arlen),   //                  .arlen
		.h2f_ARSIZE         (h2f_axi_master_arsize),  //                  .arsize
		.h2f_ARBURST        (h2f_axi_master_arburst), //                  .arburst
		.h2f_ARLOCK         (h2f_axi_master_arlock),  //                  .arlock
		.h2f_ARCACHE        (h2f_axi_master_arcache), //                  .arcache
		.h2f_ARPROT         (h2f_axi_master_arprot),  //                  .arprot
		.h2f_ARVALID        (h2f_axi_master_arvalid), //                  .arvalid
		.h2f_ARREADY        (h2f_axi_master_arready), //                  .arready
		.h2f_RID            (h2f_axi_master_rid),     //                  .rid
		.h2f_RDATA          (h2f_axi_master_rdata),   //                  .rdata
		.h2f_RRESP          (h2f_axi_master_rresp),   //                  .rresp
		.h2f_RLAST          (h2f_axi_master_rlast),   //                  .rlast
		.h2f_RVALID         (h2f_axi_master_rvalid),  //                  .rvalid
		.h2f_RREADY         (h2f_axi_master_rready),  //                  .rready
		.f2h_axi_clk        (clk_clk),                //     f2h_axi_clock.clk
		.f2h_AWID           (),                       //     f2h_axi_slave.awid
		.f2h_AWADDR         (),                       //                  .awaddr
		.f2h_AWLEN          (),                       //                  .awlen
		.f2h_AWSIZE         (),                       //                  .awsize
		.f2h_AWBURST        (),                       //                  .awburst
		.f2h_AWLOCK         (),                       //                  .awlock
		.f2h_AWCACHE        (),                       //                  .awcache
		.f2h_AWPROT         (),                       //                  .awprot
		.f2h_AWVALID        (),                       //                  .awvalid
		.f2h_AWREADY        (),                       //                  .awready
		.f2h_AWUSER         (),                       //                  .awuser
		.f2h_WID            (),                       //                  .wid
		.f2h_WDATA          (),                       //                  .wdata
		.f2h_WSTRB          (),                       //                  .wstrb
		.f2h_WLAST          (),                       //                  .wlast
		.f2h_WVALID         (),                       //                  .wvalid
		.f2h_WREADY         (),                       //                  .wready
		.f2h_BID            (),                       //                  .bid
		.f2h_BRESP          (),                       //                  .bresp
		.f2h_BVALID         (),                       //                  .bvalid
		.f2h_BREADY         (),                       //                  .bready
		.f2h_ARID           (),                       //                  .arid
		.f2h_ARADDR         (),                       //                  .araddr
		.f2h_ARLEN          (),                       //                  .arlen
		.f2h_ARSIZE         (),                       //                  .arsize
		.f2h_ARBURST        (),                       //                  .arburst
		.f2h_ARLOCK         (),                       //                  .arlock
		.f2h_ARCACHE        (),                       //                  .arcache
		.f2h_ARPROT         (),                       //                  .arprot
		.f2h_ARVALID        (),                       //                  .arvalid
		.f2h_ARREADY        (),                       //                  .arready
		.f2h_ARUSER         (),                       //                  .aruser
		.f2h_RID            (),                       //                  .rid
		.f2h_RDATA          (),                       //                  .rdata
		.f2h_RRESP          (),                       //                  .rresp
		.f2h_RLAST          (),                       //                  .rlast
		.f2h_RVALID         (),                       //                  .rvalid
		.f2h_RREADY         (),                       //                  .rready
		.h2f_lw_axi_clk     (clk_clk),                //  h2f_lw_axi_clock.clk
		.h2f_lw_AWID        (),                       // h2f_lw_axi_master.awid
		.h2f_lw_AWADDR      (),                       //                  .awaddr
		.h2f_lw_AWLEN       (),                       //                  .awlen
		.h2f_lw_AWSIZE      (),                       //                  .awsize
		.h2f_lw_AWBURST     (),                       //                  .awburst
		.h2f_lw_AWLOCK      (),                       //                  .awlock
		.h2f_lw_AWCACHE     (),                       //                  .awcache
		.h2f_lw_AWPROT      (),                       //                  .awprot
		.h2f_lw_AWVALID     (),                       //                  .awvalid
		.h2f_lw_AWREADY     (),                       //                  .awready
		.h2f_lw_WID         (),                       //                  .wid
		.h2f_lw_WDATA       (),                       //                  .wdata
		.h2f_lw_WSTRB       (),                       //                  .wstrb
		.h2f_lw_WLAST       (),                       //                  .wlast
		.h2f_lw_WVALID      (),                       //                  .wvalid
		.h2f_lw_WREADY      (),                       //                  .wready
		.h2f_lw_BID         (),                       //                  .bid
		.h2f_lw_BRESP       (),                       //                  .bresp
		.h2f_lw_BVALID      (),                       //                  .bvalid
		.h2f_lw_BREADY      (),                       //                  .bready
		.h2f_lw_ARID        (),                       //                  .arid
		.h2f_lw_ARADDR      (),                       //                  .araddr
		.h2f_lw_ARLEN       (),                       //                  .arlen
		.h2f_lw_ARSIZE      (),                       //                  .arsize
		.h2f_lw_ARBURST     (),                       //                  .arburst
		.h2f_lw_ARLOCK      (),                       //                  .arlock
		.h2f_lw_ARCACHE     (),                       //                  .arcache
		.h2f_lw_ARPROT      (),                       //                  .arprot
		.h2f_lw_ARVALID     (),                       //                  .arvalid
		.h2f_lw_ARREADY     (),                       //                  .arready
		.h2f_lw_RID         (),                       //                  .rid
		.h2f_lw_RDATA       (),                       //                  .rdata
		.h2f_lw_RRESP       (),                       //                  .rresp
		.h2f_lw_RLAST       (),                       //                  .rlast
		.h2f_lw_RVALID      (),                       //                  .rvalid
		.h2f_lw_RREADY      ()                        //                  .rready
	);

endmodule
