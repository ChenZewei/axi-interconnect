library verilog;
use verilog.vl_types.all;
entity axi_interface is
end axi_interface;
